package enums;

   typedef enum
   {
       IDLE,
       SHIFT_1,
       SHIFT_2,
       SHIFT_3,
       HOLDING
   } state_t;

endpackage

